`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    12:51:20 04/20/2019 
// Design Name: 
// Module Name:    id_ex_reg 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module id_ex_reg(
	 input clk,
    input rst,
    input data_input,
    input control_data_input,
    output data_output,
    output control_data_output
    );


endmodule
